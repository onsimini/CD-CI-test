module top(
    input   wire    i_switch,
    output  wire    o_led
);

    assign  o_led = i_switch;

endmodule
